-- alarm 闹铃模块

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY alarm IS
    PORT (
		  SET_HOUR10: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  SET_HOUR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  SET_MIN10: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  SET_MIN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  HOUR10: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  HOUR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  MIN10: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  MIN: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  SEC10: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  SEC: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  SPEAKER: OUT STD_LOGIC
		 );
END alarm;
ARCHITECTURE behavioral OF alarm IS	
	BEGIN
		clock_alarm:PROCESS(SET_HOUR10, SET_HOUR, SET_MIN10, SET_MIN,
		HOUR10, HOUR, MIN10, MIN, SEC10, SEC)
		BEGIN
			IF SEC10 = "0001" THEN
				SPEAKER <= '0';
			ELSIF SEC10 = "0100" THEN
				SPEAKER <= '0';
			ELSIF SEC = "0100" THEN
				SPEAKER <= '0';
			ELSIF MIN10 = "0101" AND MIN = "1001" AND SEC10 = "0101" AND SEC = "0101" THEN
				SPEAKER <= '1';
			ELSIF MIN10 = "0101" AND MIN = "1001" AND SEC10 = "0101" AND SEC = "0111" THEN
				SPEAKER <= '1';
			ELSIF MIN10 = "0101" AND MIN = "1001" AND SEC10 = "0101" AND SEC = "1001" THEN
				SPEAKER <= '1';
			ELSIF HOUR10 = SET_HOUR10 AND HOUR = SET_HOUR AND MIN10 = SET_MIN10 AND MIN = SET_MIN AND SEC10 = "0000" THEN
				SPEAKER <= '1';
			ELSE SPEAKER <= '0';
			END IF;
		END PROCESS;
END behavioral;